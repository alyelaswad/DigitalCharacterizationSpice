CMOS Inverter Analysis
.include MOSFET_models_0p5_0p18-1.inc
VIN 1 0 PULSE(3.3 0 0 0.1n 0.1n 10n 20n)  ; Pulse input with rise and fall times of 0.1n and period 20n
VVDD 3 0 DC 3.3
M1 2 1 0 0 NMOS0P5 [w=1.25u l=0.5u As=1.875p Ad=1.875p ps=5.5u pd=5.5u]
M2 2 1 3 3 PMOS0P5 [w=1.25u l=0.5u As=1.875p Ad=1.875p ps=5.5u pd=5.5u]
RL 2 4 1k
CL 4 0 0.5p
.tran 1n 20n; Transient analysis for one period of the input (20ns)
.END
